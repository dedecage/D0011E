library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Programmemory is
    Port ( Address:in std_logic_vector(31 downto 0);
           Instruction: out std_logic_vector(31 downto 0));
end Programmemory;

architecture behav of Programmemory is
begin

with address select
  instruction <="00100000001000001111111111111000" when X"00000000",  --addi r0,r1,-8 | r0 = -8 | -8
                "00100000010000010000000000000011" when X"00000004",  --addi r1,r2,3 | r1 = 3 | 3
		        "00000000000000010001000000100000" when X"00000008",  --add r2,r0,r1 | r2 = -5 | 3
                "00000000001000000001100000100010" when X"0000000c",  --sub r3,r1,r0 | r3 = 11 | 3
		        "00000000010000110010000000101010" when X"00000010",  --slt r4,r2,r3 | r4 = 1 | 0
		        "00101000010001001111111111110111" when X"00000014",  --slti r4,r2,-9 | r4 = 0 | 0
		        "00000000010000110010000000101010" when X"00000018",  --slt r4,r2,r3 | r4 = 1 | 0
		        "00000000100001100010100000100101" when X"0000001c",  --or  r5,r4,r6 | r5 = 1 | 0
		        "00000000101000010011000000100100" when X"00000020",  --and r6,r5,r1 | r6 = 1 | 0
		        "10101100111000100000000000000000" when X"00000024",   --sw r2, 0(r7)  | r2 = (0+r7)
                "10001100111010000000000000000000" when X"00000028",   --lw r8, 0(r7)  | r8 = (0+r8)
                "10101101001000110000000000000100" when X"0000002c",   --sw r3, 4(r9)  | r3 = (4+r9)
                "10001101010010010000000000000100" when X"00000030",   --lw r9, 4(r10) | r9 = (4+r10)
                "11111100001000000000000000000001" when others;
                
-- TEST N = 12, D = 5              
--instruction <=  "00100000000000100000000000000000" when X"00000000", --addi $r2, $r0, 0 -- Q = 0  
--                "00100000000001000000000000001100" when X"00000004", --addi $r4, $r0, 0x000c, N = 12
--                "00100000000001010000000000000101" when X"00000008", --addi $r5, $r0, 0x0005, D = 5
--                "00100000100000110000000000000000" when X"0000000c", --addi $r3, $r4, 0x0000, R = N
--                "00100000000001100000000000000001" when X"00000010", --addi $r6, r0, 1
--                "00000000011001010011100000101010" when X"00000014", --slt $r7, $r3, $r5
--                "00010000110001110000000000000011" when X"00000018", --beq $r6, $r7, 3
--                "00100000010000100000000000000001" when X"0000001c", --addi $r2, $r2, 1
--                "00000000011001010001100000100010" when X"00000020", --sub $r3, $r3, $r5
--                "00001000000000000000000000000100" when X"00000024", --j 4
--                "10101100000000100000000000000010" when X"00000028", --sw $r2, 2($r0)
--                "10101100000000110000000000000011" when X"0000002c", --sw $r3, 3($r0)
                
       
-- TEST N = 12, D = 12 
--instruction <=  "00100000000000100000000000000000" when X"00000000", --addi $r2, $r0, 0 -- Q = 0
--                "00100000000001000000000000001100" when X"00000004", --addi $r4, $r0, 0x000c, N = 12
--                "00100000000001010000000000001100" when X"00000008", --addi $r5, $r0, 0x0005, D = 12
--                "00100000100000110000000000000000" when X"0000000c", --addi $r3, $r4, 0x0000, R = N
--                "00100000000001100000000000000001" when X"00000010", --addi $r6, r0, 1
--                "00000000011001010011100000101010" when X"00000014", --slt $r7, $r3, $r5
--                "00010000110001110000000000000011" when X"00000018", --beq $r6, $r7, 3
--                "00100000010000100000000000000001" when X"0000001c", --addi $r2, $r2, 1
--                "00000000011001010001100000100010" when X"00000020", --sub $r3, $r3, $r5
--                "00001000000000000000000000000100" when X"00000024", --j 4
--                "10101100000000100000000000000010" when X"00000028", --sw $r2, 2($r0)
--                "10101100000000110000000000000011" when X"0000002c", --sw $r3, 3($r0)
   
---- TEST N = 5, D = 12
--   instruction <=  "00100000000000100000000000000000" when X"00000000", --addi $r2, $r0, 0 -- Q = 0
--                   "00100000000001000000000000000101" when X"00000004", --addi $r4, $r0, 0x0005, N = 5
--                   "00100000000001010000000000001100" when X"00000008", --addi $r5, $r0, 0x0005, D = 12
--                   "00100000100000110000000000000000" when X"0000000c", --addi $r3, $r4, 0x0000, R = N
--                   "00100000000001100000000000000001" when X"00000010", --addi $r6, r0, 1
--                   "00000000011001010011100000101010" when X"00000014", --slt $r7, $r3, $r5
--                   "00010000110001110000000000000011" when X"00000018", --beq $r6, $r7, 3
--                   "00100000010000100000000000000001" when X"0000001c", --addi $r2, $r2, 1
--                   "00000000011001010001100000100010" when X"00000020", --sub $r3, $r3, $r5
--                   "00001000000000000000000000000100" when X"00000024", --j 4
--                   "10101100000000100000000000000010" when X"00000028", --sw $r2, 2($r0)
--                   "10101100000000110000000000000011" when X"0000002c", --sw $r3, 3($r0)

end behav;

